// Sample 5.27 Good transactions creator task with ref on handle

function void create(ref Transaction tr);
	///...
	
endfunction : create