// Sample 6.36 $urandom_range usage

a = $urandom_range(3,10);			// Pick a value from 3 to 10
a = $urandom_range(10,3);			// Pick a value from 3 to 10
b = $urandom_range(5);				// Pick a value from 0 to 5
