// Sample 5.2 Class in a package


package abc;
	class Transaction;
		//Class body
	endclass : Transaction
endpackage : abc