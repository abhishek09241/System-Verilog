// Sample 5.17 Static method displays static variable

class Transaction;
	static Config cfg;				// A handle with static storage