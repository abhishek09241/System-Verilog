// Sample 5.3 Shows hot to import a package into a program


program automatic test;
	import abc::*;
	Transaction tr;			// Declare a handle  and value of (tr is null)
	tr = new();				// Allocate a Transaction object


	// Test code
	
endprogram