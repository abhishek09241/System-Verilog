// Sample 8.40 Transactor class with static print class

class Xactor
	task run();
		Print::error("NYI","This Xactor is not yet implemented");
	endtask : run

endclass: Xactor